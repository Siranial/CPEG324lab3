library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity comparator is
    Port (  A,B : in STD_LOGIC_VECTOR (7 downto 0);
            S : in STD_LOGIC;
            Y : out STD_LOGIC_vector (7 downto 0));
end comparator;

architecture Behavioral of comparator is

begin

    -- Logic

end Behavioral;