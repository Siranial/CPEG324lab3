library ieee;
use ieee.std_logic_1164.all;

entity alu is
    Port (  
    );
end alu;

architecture behavioral of alu is

    -- Component Instantiation

    begin

        -- Logic

end behavioral;